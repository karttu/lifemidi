/* lifemidi.v   --   Copyright (C) 2005-2012, Antti Karttunen.

   A module for Spartan-3 Starter Board, which iterates Conway's Life on
   Mefisto 8x8 chess board, while at the same time iterating permutations
   of eight elements, and producing MIDI-music based on those inputs.

   For interesting patterns of dynamics, check http://oeis.org/A179409
   and http://oeis.org/A179412 especially the latter.

   Unless otherwise mentioned, all Verilog-modules in this code tree are
   Copyright (C) 2010-2012 Antti Karttunen, subject to the terms of the GPL v2.
   See the file COPYING for more information.  Contact the author for further
   developments at the address <his-firstname>.<his-surname>@gmail.com


   Changes, some of them:

   An early version from January 29 2010 adds the population & generation counts
   (the former is shown in two rightmost 7-seg led digits, while the leftmost
    8 bits of the latter are shown as binary in the leds LD0--LD7.)

   Also as a novelty we have non-single-stepped operation. Switches 5-0 determine the
   running speed, from 1.514 Hz to 95.4 Hz. If they are all in 0-position,
   then we run in single-step mode.

   Version March 24 2010 added MIDI-output. Now the pauses are four times slower,
   so that there's enough time to play all eight notes between each generation.

   Version March 25 2010 with external SYNC -input.
	
   First somehow working version (of MIDI), 10:50 am Mar 26 2010.
   Turning notes off works now as expected.

   The population count still shows the _previous_ generation.
    
   Now the demanded feature: the ext sync divider.
   Its settings work in funny way, not all push buttons completely independent.
   (This version, Mar 26 2010, 1:25 pm).

   New version, April 06 & 07 2010:

   Switch 0 determines how the the MIDI-notes are turned off:

    When in high position (1), the notes are not turned off,
                               until before the next round,
                               they might be turned off,
                               if that row is at that time all zeroes.
    When in low position (0),  the notes are turned off before
                               the next one is turned on.

   Switch 1 determines how the velocity value for each note
   is contructed.

    When in low position (0), it's copied directly from the seven
                              least significant bits of each row.

    When in high position (1), it's just the number of alive cells
                               on that row * 16 - 1 (if not zero), to get values
                               (0, 16, 32, 48, 64, 80, 96, 112, 128)
                               (0, 15, 31, 47, 63, 79, 95, 111, 127).


    Version 07 April with permuting of the scale.
    (Bug: zero-rows don't generate zero-velocity in alive-cell-count mode.)

    Development continued on October 6th 2012.
    The name of design and the top-module changed to lifemidi.
    Added Digitel-2000 16x7 seg led display. (For showing the factorial
    expansion and the associated permutation.)
 
    2012-10-08: Merged with the most important additions of the
    version 24 April 2010, where the above zero-rows bug was fixed, and also
    with the detection of stable/oscillating-period-2 patterns,
    whence a new Life-pattern is copied from the permutation when
    such a stagnated situation has been detected.

    2012-10-10: Added the initialization of factorial expansion/permutation
                with Ericsson rotary dialer.

    2012-10-20: Added a new argument invert_sync_in to syncdivider module.
                Testing the dialer-syncing.

 */

module lifemidi(input CLK, // 50Mhz internal clock of Spartan-3 XC200 FPGA.
                input [3:0] PB_IN, // Push-buttons in Spartan-3 Starter Board
                input DIN_SYNC_IN, // External sync coming with "MIDI-cable"
//                                    (i.e. 5-pin DIN) thru optoisolater board.
                input [7:0] SW_IN, // Switches in Spartan-3 Starter Board.

                input dialer_in_rest, // HI if dialer is in its rest-position.
//                             Thru "sidewing" at User B1 Expansion Connector.
                input dialer_pulses,  // Pulses generated by dialer.

// The next three go through the optoisolator-board, and are all optoisolated:
                input [7:0] BCOL_IN,  // Which reed-relays are closed on the
// currently sampled (multiplexed) row of Mefisto-matrix?
                output [7:0] BCOL_OUT, // Show these leds on the currently
// multiplexed row of Mefisto-matrix.
                output [7:0] BROW,    // For multiplexing the rows of Mefisto
// LED & Reed-relay matrix. Used as rotating one-hot shift-register.

                output [7:0] LED_OUT, // Eight leds on Spartan-3 Starter Board.
                output [7:0] SEG_OUT, // The segments of four LED-digits on SP3
                output [3:0] DIGIT_OUT, // Which digit to show? Rotate one-cold
//                                         (They seem to be inverted common anodes)

                output MIDIOUT,       // Where the midi-notes are sent. This
// is via a transistor located on optoisolater-board. (This signal is not
// optoisolated on our end. The transistor's emitter is connected to the
// grounds of both 3,3V and 5V side of the OI-board, so the sides are
// not anymore galvanically separated.)

                output [7:0] extseg_out, // The segments of 16 LED-digits on
// Digitel-2000 display. Thru User B1 Extension Port side-wing.
                output [15:0] extdigit_out // The common cathodes for eight
// segments of each of the digits. Use multiplexed one-cold rotating shift-reg.
               );

reg [15:0] main_cycle_ctr = 16'b0000000000000001;
// wire RST = PB_IN[3];


reg [7:0] BOARD_ROW [7:0];
reg [7:0] PREV1_BOARD_ROW [7:0];
reg [7:0] PREV2_BOARD_ROW [7:0];

wire [7:0] PIECES_ROW [7:0];

// If we xor the current board with the situation two generations ago,
// and the result is zero, then we have either fallen into a stable
// pattern (including dead ones) or one oscillating with period 2:
wire has_stagnated = ~(|(PREV2_BOARD_ROW[0]^BOARD_ROW[0])
                     | |(PREV2_BOARD_ROW[1]^BOARD_ROW[1])
                     | |(PREV2_BOARD_ROW[2]^BOARD_ROW[2])
                     | |(PREV2_BOARD_ROW[3]^BOARD_ROW[3])
                     | |(PREV2_BOARD_ROW[4]^BOARD_ROW[4])
                     | |(PREV2_BOARD_ROW[5]^BOARD_ROW[5])
                     | |(PREV2_BOARD_ROW[6]^BOARD_ROW[6])
                     | |(PREV2_BOARD_ROW[7]^BOARD_ROW[7])
                     );

reg [3:0] rs[7:0]; // The row sums.
reg [6:0] rv[7:0]; // The row velocities, computed from the sums.

reg [6:0] popula = 7'b0000000; // Population count. From 0 to 64.
reg [6:0] old_popula = 7'b1111111; // Its contents in the prev cycle.
reg [15:0] this_generation = 0;

// wire [2:0] shrow = {SW_IN[2],SW_IN[1],SW_IN[0]};

wire input_mode = SW_IN[7];

wire notes_turned_off     = ~SW_IN[0];
wire note_velocity_summed = SW_IN[1];


// wire [5:0] selected_speed = SW_IN[5:0];
// wire [5:0] selected_speed = {SW_IN[6:3]}; // Our switch 2 has jammed.
wire [3:0] selected_speed = {SW_IN[6:3]};

// Compute the pause period from the speed selection switches:
function [24:0] get_pp;
  input [3:0] ss; // Speed switches 3:0.~ss[3],~ss[4],~ss[5]
  get_pp = ({~ss[0],~ss[1],~ss[2],~ss[3],1'b0,1'b0}+6'b000001) << 19;
endfunction


function fredkin;
  input n;
  input s;
  input w;
  input e;
  fredkin = (n^s^w^e);
endfunction


// The cell will be alife if it has either 3 neighbours
// or if it has 2 neighbours and it itself is alive.
function life;
  input c;
  input n;
  input ne;
  input s;
  input se;
  input w;
  input sw;
  input e;
  input nw;
//life = (4'b0011 == ((n+ne+e+se+s+sw+w+nw)|c));
  life = (4'b0011 == (({3'b000,n}+{3'b000,ne}+{3'b000,s}+{3'b000,se}+{3'b000,w}+{3'b000,sw}+{3'b000,e}+{3'b000,nw})|{3'b000,c}));
endfunction

function [3:0] c8b;
  input [7:0] b;
  c8b = ({3'b000,b[7]}+{3'b000,b[6]}+{3'b000,b[5]}+{3'b000,b[4]}+{3'b000,b[3]}+{3'b000,b[2]}+{3'b000,b[1]}+{3'b000,b[0]});
endfunction

function [30:0] rol31bits;
  input [30:0] b;
  rol31bits = {b[29],b[28],b[27],b[26],b[25],b[24],b[23],b[22],b[21],b[20],
                b[19],b[18],b[17],b[16],b[15],b[14],b[13],b[22],b[11],b[10],
                b[9],b[8],b[7],b[6],b[5],b[4],b[3],b[2],b[1],b[0],b[30]};
endfunction

// This doesn't rotate, but just shifts left, and fills bit-zero with zero.
function [30:0] shl31bits;
  input [30:0] b;
  shl31bits = {b[29],b[28],b[27],b[26],b[25],b[24],b[23],b[22],b[21],b[20],
                b[19],b[18],b[17],b[16],b[15],b[14],b[13],b[22],b[11],b[10],
                b[9],b[8],b[7],b[6],b[5],b[4],b[3],b[2],b[1],b[0],1'b0};
endfunction


mefi8x8a BOARD_IO(.CLK(CLK),
                  .BCOL_IN(BCOL_IN),
                  .BCOL_OUT(BCOL_OUT),
                  .BROW(BROW),
                  .LEDS2LIT0(BOARD_ROW[0]),
                  .LEDS2LIT1(BOARD_ROW[1]),
                  .LEDS2LIT2(BOARD_ROW[2]),
                  .LEDS2LIT3(BOARD_ROW[3]),
                  .LEDS2LIT4(BOARD_ROW[4]),
                  .LEDS2LIT5(BOARD_ROW[5]),
                  .LEDS2LIT6(BOARD_ROW[6]),
                  .LEDS2LIT7(BOARD_ROW[7]),
                  .PIECES0(PIECES_ROW[0]),
                  .PIECES1(PIECES_ROW[1]),
                  .PIECES2(PIECES_ROW[2]),
                  .PIECES3(PIECES_ROW[3]),
                  .PIECES4(PIECES_ROW[4]),
                  .PIECES5(PIECES_ROW[5]),
                  .PIECES6(PIECES_ROW[6]),
                  .PIECES7(PIECES_ROW[7])
                 );


wire use_dialer_for_beat = SW_IN[2];
wire dialer_debounced_pulses;

wire SYNC_IN = (use_dialer_for_beat ? dialer_debounced_pulses : DIN_SYNC_IN);

reg SYNC_IN_S = 0;
reg SYNC_IN_S_PREV = 0;

wire pb0_next; // State of the debounced push button for incrementing.
reg pb0_next_prev = 0; // is saved here also.

wire pb1_next; // State of the debounced push button for incrementing.
reg pb1_next_prev = 0; // is saved here also.

wire pb2_next; // State of the debounced push button for incrementing.
reg pb2_next_prev = 0; // is saved here also.


wire pb0_pressed = (pb0_next && ~pb0_next_prev);
wire pb1_pressed = (pb1_next && ~pb1_next_prev);
wire pb2_pressed = (pb2_next && ~pb2_next_prev);

debounced_button DBB0(CLK,PB_IN[0],pb0_next);
debounced_button DBB1(CLK,PB_IN[1],pb1_next);
debounced_button DBB2(CLK,PB_IN[2],pb2_next);

wire sync_invert_sync_in;


// wire ext_sync_raised = ((SYNC_IN_S & (SYNC_IN_S!=SYNC_IN_S_PREV))| pb0_pressed);
wire ext_sync_changed = (pb0_pressed|((SYNC_IN_S ^ sync_invert_sync_in) & (SYNC_IN_S!=SYNC_IN_S_PREV)));

wire divided_sync;
// wire divided_sync = ext_sync_raised;

wire [3:0] sync_divby;
wire [3:0] sync_sel_offset;

syncdivider SYNCDIV(.CLK(CLK),
                    .sync_in(ext_sync_changed),
                    .sync_out(divided_sync),
                    .pb_divby(pb2_pressed),
                    .pb_offset(pb1_pressed),
                    .divby(sync_divby),
                    .sel_offset(sync_sel_offset),
                    .invert_sync_in(sync_invert_sync_in)
                   );

// 2^19 * 20ns = 524288 * 20 ns = 0.0105 sec = 10.5 ms. (95.4 Hz)
// 63 * 10.5 ms = 0.66 sec (1.51 Hz)
// reg [24:0] pause_counter = 25'b0000000000000000000000000;

// 2^21 * 20ns = 2097152 * 20 ns = 0.0419 sec = 42 ms. (23.8 Hz)
// 63 * 42 ms = 2.646 sec (0.38 Hz)

// 2^22 * 20ns = 4194304 * 20 ns = 0.083886 sec = 84 ms. (11.9 Hz)
// 63 * 84 ms = 5.285 sec (0.189 Hz) / 8 = 0.66060288 sec.

reg [24:0] pause_counter = 25'b0000000000000000000000000;

// We proceed to play the next midi-note when either
// a) the user has selected non-zero pause-period (i.e. not single-step)
//    and the pause period has just completed (it's all zeros),
// or
// b) single_step button has been pressed:
 
// wire sync_signal = ((|selected_speed & ~|pause_counter) | ext_sync_raised);
wire sync_signal = ((|selected_speed & ~|pause_counter) | divided_sync);

reg [2:0] row_index = 3'b000;
reg [2:0] next_row_index = 3'b000;


function [7:0] OCT2HOTCODE;
  input [2:0] OCT;

  begin
    case (OCT)
      3'b001  : OCT2HOTCODE = 8'b00000010;	//1
      3'b010  : OCT2HOTCODE = 8'b00000100;	//2
      3'b011  : OCT2HOTCODE = 8'b00001000;	//3
      3'b100  : OCT2HOTCODE = 8'b00010000;	//4
      3'b101  : OCT2HOTCODE = 8'b00100000;	//5
      3'b110  : OCT2HOTCODE = 8'b01000000;	//6
      3'b111  : OCT2HOTCODE = 8'b10000000;	//7
      default : OCT2HOTCODE = 8'b00000001;	//0
    endcase
  end
endfunction


function [6:0] OCT2NBITS_FROM_RIGHT;
  input [2:0] OCT;

  begin
    case (OCT)
      3'b001  : OCT2NBITS_FROM_RIGHT = 7'b0000001;	//1
      3'b010  : OCT2NBITS_FROM_RIGHT = 7'b0000011;	//2
      3'b011  : OCT2NBITS_FROM_RIGHT = 7'b0000111;	//3
      3'b100  : OCT2NBITS_FROM_RIGHT = 7'b0001111;	//4
      3'b101  : OCT2NBITS_FROM_RIGHT = 7'b0011111;	//5
      3'b110  : OCT2NBITS_FROM_RIGHT = 7'b0111111;	//6
      3'b111  : OCT2NBITS_FROM_RIGHT = 7'b1111111;	//7
      default : OCT2NBITS_FROM_RIGHT = 7'b0000000;	//0
    endcase
  end
endfunction


////////   MIDI OUTPUT   /////////

// int scale_pentatonic_minor[] = { 0, 3, 5, 7, 10, 12, 15, 17 };

function [7:0] pentatonic_minor_C4;
  input [2:0] relnote;
  begin
    case (relnote)
      3'd0 : pentatonic_minor_C4 = 8'd60 + 8'd17;
      3'd1 : pentatonic_minor_C4 = 8'd60 + 8'd15;
      3'd2 : pentatonic_minor_C4 = 8'd60 + 8'd12;
      3'd3 : pentatonic_minor_C4 = 8'd60 + 8'd10;
      3'd4 : pentatonic_minor_C4 = 8'd60 + 8'd7;
      3'd5 : pentatonic_minor_C4 = 8'd60 + 8'd5;
      3'd6 : pentatonic_minor_C4 = 8'd60 + 8'd3;
      default : pentatonic_minor_C4 = 8'd60 + 8'd0;
    endcase
  end
endfunction

wire [2:0] midibeat = row_index;


parameter initial31onehot = 31'b0000000000000000000000000000001;

// This is one hot register:
reg [30:0] syncdelay = initial31onehot;
wire [30:0] nextsyncdelay = (sync_signal ? initial31onehot : (syncdelay << 1));
 

// We have to take care, that when sync_signal comes,
// we do these things in order:
//  a) Turn off the previous note, for the current row_index
//  b) Increment the row index, after some safe delay from (a).
//    c) If the new row index is zero, i.e. we have scanned all
//       eight rows/pitches, compute the next Life-generation.
//    d) permute the scale.
//  f) Turn on the next note, for the current incremented row_index,
//       after some safe delay from (b), (c) and (d).

parameter time_one_after_beat    = 0;
parameter time2turn_off_prevnote = 0;
parameter time2comp_next_gen     = 6;
parameter time2comp_next_perm    = 7;
parameter time2sum_the_rows      = 8;
parameter time2comp_velocities   = 9;
parameter time2inc_to_next_row   = 10;
parameter time2turn_on_nextnote  = 15;
parameter time2showpopcnt        = 30;


wire show_pop_count = ((syncdelay[time2showpopcnt])
                       | (input_mode && (popula != old_popula))
                       | pb0_pressed | pb1_pressed | pb2_pressed);



wire comp_next_gen = (~|next_row_index & (syncdelay[time2comp_next_gen]));

wire [24:0] next_pause_counter
  = ((input_mode|syncdelay[time_one_after_beat]) ? get_pp(selected_speed)
                                                  : (pause_counter-1));


// Turn the prev note off immediately at sync rising edge.
wire midinoteoff = (notes_turned_off & syncdelay[time2turn_off_prevnote]);
wire midinoteon  = syncdelay[time2turn_on_nextnote];
wire midisendtriplet = (midinoteoff | midinoteon);


wire [2:0] op [7:0]; // From perm8eng.

wire [7:0] midinote = pentatonic_minor_C4(op[midibeat]);

// assign LED_OUT = this_generation[7:0];
assign LED_OUT[2:0] = row_index;
assign LED_OUT[6:3] = selected_speed[3:0]; // Just for debugging

assign LED_OUT[7] = SYNC_IN; // sync_signal; // Testing.

wire [7:0] midivelocity = (midinoteoff ? 0 : {1'b0,rv[midibeat]});

// wire [7:0] midivelocity = (midinoteoff ? 0 : {1'b0,rv[midibeat]});

//                            : {1'b0,BOARD_ROW[midibeat][6:0]});
//                            : (0==midibeat) ? {1'b0,BOARD_ROW[0][6:0]}
//                            : (1==midibeat) ? {1'b0,BOARD_ROW[1][6:0]}
//                            : (2==midibeat) ? {1'b0,BOARD_ROW[2][6:0]}
//                            : (3==midibeat) ? {1'b0,BOARD_ROW[3][6:0]}
//                            : (4==midibeat) ? {1'b0,BOARD_ROW[4][6:0]}
//                            : (5==midibeat) ? {1'b0,BOARD_ROW[5][6:0]}
//                            : (6==midibeat) ? {1'b0,BOARD_ROW[6][6:0]}
//                            : {1'b0,BOARD_ROW[7][6:0]}
//                          );


midiout3bytes MIDINoteOnOff(.CLK(CLK),
                            .RST(PB_IN[3]), // User reset for MIDI-Uart.
                            .ibyte1(8'h90),
                            .ibyte2(midinote),
                            .ibyte3(midivelocity),
                            .sendthem(midisendtriplet),
                            .MIDIOUT(MIDIOUT)
                           );

///////// PERMUTATION ENGINE & ITS INITIALIZATION WITH DIALER /////////

reg prev_all_digits_dialed = 1'b0;
// Raise it up for just one cycle:
wire all_digits_dialed;
wire [2:0] n_digits_dialed;

wire all_digits_just_dialed = (~prev_all_digits_dialed & all_digits_dialed);

wire synced_dialer_in_rest;

syncinp SYNC_RESTSIGNAL(CLK,dialer_in_rest,synced_dialer_in_rest);

// As long as dialer is not in rest or not all digits have been dialed
wire is_dialing = (~synced_dialer_in_rest) | ~all_digits_dialed;
// De Morgan: ~(dialer_in_rest & all_digits_dialed);


wire       of1;
wire [1:0] of2;
wire [1:0] of3;
wire [2:0] of4;
wire [2:0] of5;
wire [2:0] of6;
wire [2:0] of7;

// For user-dialed 7-digit factorial expansion, 0000000 .. 7654321

wire dialed_f1;         // 0-1
wire [1:0]  dialed_f2;  // 0-2
wire [1:0]  dialed_f3;  // 0-3
wire [2:0]  dialed_f4;  // 0-4
wire [2:0]  dialed_f5;  // 0-5
wire [2:0]  dialed_f6;  // 0-6
wire [2:0]  dialed_f7;  // 0-7

wire show_f1 = (is_dialing ? dialed_f1 : of1);
wire [1:0] show_f2 = (is_dialing ? dialed_f2 : of2);
wire [1:0] show_f3 = (is_dialing ? dialed_f3 : of3);
wire [2:0] show_f4 = (is_dialing ? dialed_f4 : of4);
wire [2:0] show_f5 = (is_dialing ? dialed_f5 : of5);
wire [2:0] show_f6 = (is_dialing ? dialed_f6 : of6);
wire [2:0] show_f7 = (is_dialing ? dialed_f7 : of7);


   
wire permreset = (input_mode | all_digits_just_dialed);

wire next_perm = (~|next_row_index & (syncdelay[time2comp_next_perm]));

wire [2:0] zero_triplet = 3'b000;

wire inf1 = (all_digits_dialed ? dialed_f1 : zero_triplet);
wire [1:0] inf2 = (all_digits_dialed ? dialed_f2 : zero_triplet);
wire [1:0] inf3 = (all_digits_dialed ? dialed_f3 : zero_triplet);
wire [2:0] inf4 = (all_digits_dialed ? dialed_f4 : zero_triplet);
wire [2:0] inf5 = (all_digits_dialed ? dialed_f5 : zero_triplet);
wire [2:0] inf6 = (all_digits_dialed ? dialed_f6 : zero_triplet);
wire [2:0] inf7 = (all_digits_dialed ? dialed_f7 : zero_triplet);


perm8eng PERMENGINE(CLK,
                    permreset,
                    next_perm,
                    inf1,inf2,inf3,inf4,inf5,inf6,inf7,
                    of1,of2,of3,of4,of5,of6,of7,
                    op[0],op[1],op[2],op[3],
                    op[4],op[5],op[6],op[7]);


dialerfe DIALER(.CLK(CLK),
                .restart(input_mode | all_digits_just_dialed),
                .dialer_in_rest(synced_dialer_in_rest),
                .dialer_pulses(dialer_pulses),
                .all_digits_have_been_dialed(all_digits_dialed),
                .num_of_digits_dialed(n_digits_dialed),
                .of1(dialed_f1),
                .of2(dialed_f2),
                .of3(dialed_f3),
                .of4(dialed_f4),
                .of5(dialed_f5),
                .of6(dialed_f6),
                .of7(dialed_f7),
                .debounced_pulses(dialer_debounced_pulses));



///////// FOUR DIGIT SPARTAN-3 DEVBOARD 7-SEG DISPLAY /////////


// shw16decb DECDISPLAY(CLK,butbuf[7],this_generation[15:0],SEG_OUT,DIGIT_OUT);
// shw16decb DECDISPLAY(CLK,show_pop_count,{9'b000000000,popula[6:0]},SEG_OUT,DIGIT_OUT);

// shw16decb DECDISPLAY(CLK,
//                     show_pop_count,
//                     (1000*sync_divby)+(100*sync_sel_offset)+popula[6:0],
//                     SEG_OUT,DIGIT_OUT);

show16withdps DECDISPLAY(CLK,
                     show_pop_count,
// /* Debug: */      ((1000*n_digits_dialed)+(100*sync_sel_offset)+popula[6:0]),
                     ((1000*sync_divby)+(100*sync_sel_offset)+popula[6:0]),
                     all_digits_dialed,sync_invert_sync_in,dialer_pulses,synced_dialer_in_rest,
//                   all_digits_dialed,is_dialing,dialer_pulses,synced_dialer_in_rest,
                     SEG_OUT,DIGIT_OUT);



digitel2000_16x7seg PERMdisplay(.CLK(CLK),
                               .extseg_out(extseg_out),
                               .extdigit_out(extdigit_out),
                               .refresh(main_cycle_ctr[15]),
                               .dig0(op[7]),
                               .dig1(op[6]),
                               .dig2(op[5]),
                               .dig3(op[4]),
                               .dig4(op[3]),
                               .dig5(op[2]),
                               .dig6(op[1]),
                               .dig7(op[0]),
                               .dig8(3'b000), // Keep it black...
                               .dig9({2'b00,show_f1}), // Not this way! (Why not? I have forgotten why!)
                               .dig10({1'b0,show_f2}),
                               .dig11({1'b0,show_f3}),
                               .dig12(show_f4),
                               .dig13(show_f5),
                               .dig14(show_f6),
                               .dig15(show_f7),
// We do ~midibeat to get reversed indexing from 7 to 0, as op[0..7]
// are now listed from left to right.
// ~OCT2HOTCODE(~midibeat) is for showing the "ambient mode". (switch 0 up).
                               .decimal_points({8'b00000000,
                                                (notes_turned_off
                                                   ? OCT2HOTCODE(~midibeat)
                                                   : ~OCT2HOTCODE(~midibeat))
                                               }),
                               .show_only_these({(is_dialing
                                      ? OCT2NBITS_FROM_RIGHT(n_digits_dialed
                                 /* A hack! */ + {2'b00,~synced_dialer_in_rest})
                                      : 7'b1111111), // XXX - Improve!
                                                9'b011111111}));

integer i; // A "compile-time" index to board rows. (for the for loop).
integer j;

always @(posedge CLK)
  begin
   main_cycle_ctr <= main_cycle_ctr+1;
// if(RST)
//  begin
//  end
// else
//  begin
      SYNC_IN_S <= ~SYNC_IN; // Avoid metastability issues with asynchronic input.
      SYNC_IN_S_PREV <= SYNC_IN_S;

      pb0_next_prev <= pb0_next;
      pb1_next_prev <= pb1_next;
      pb2_next_prev <= pb2_next;

      prev_all_digits_dialed <= all_digits_dialed;

      pause_counter <= next_pause_counter;
      syncdelay <= nextsyncdelay;
 
      if(sync_signal)
        begin
         next_row_index <= row_index+1;
        end

      if(syncdelay[time2inc_to_next_row])
        begin
         row_index <= next_row_index;
        end


      if(input_mode)
        begin // Transfer the state from input registers (reed relays)
          old_popula <= popula;

          this_generation <= 0;
          for(i=0; i<8; i=i+1) BOARD_ROW[i] <= PIECES_ROW[i];
          for(i=0; i<8; i=i+1) PREV1_BOARD_ROW[i] <= 8'b11111111;
          for(i=0; i<8; i=i+1) PREV2_BOARD_ROW[i] <= 8'b11111111;
        end
      else if(comp_next_gen)
        begin
          old_popula <= popula;
          // Sum the population total from the current state.
          popula <= {3'b000,c8b(BOARD_ROW[0])}
                  + {3'b000,c8b(BOARD_ROW[1])}
                  + {3'b000,c8b(BOARD_ROW[2])}
                  + {3'b000,c8b(BOARD_ROW[3])}
                  + {3'b000,c8b(BOARD_ROW[4])}
                  + {3'b000,c8b(BOARD_ROW[5])}
                  + {3'b000,c8b(BOARD_ROW[6])}
                  + {3'b000,c8b(BOARD_ROW[7])};

          for(i=0; i<8; i=i+1)
           begin
            PREV2_BOARD_ROW[i] <= PREV1_BOARD_ROW[i];
            PREV1_BOARD_ROW[i] <= BOARD_ROW[i];
           end

          if(has_stagnated) // Get the new pattern from permutation:
           begin
            for(i=0; i<8; i=i+1) BOARD_ROW[i] <= {2'b00,op[i],3'b000};
           end
          else // Otherwise, compute the next Life-generation as usual:
           begin
            for(i=0; i<8; i=i+1)
             for(j=0; j<8; j=j+1)
                BOARD_ROW[i][j] <= life(BOARD_ROW[i][j], // The cell itself.
                                        BOARD_ROW[i][(7==j ? 0 : j+1)], // n
                                        BOARD_ROW[(7==i ? 0 : i+1)][(7==j ? 0 : j+1)], // ne
                                        BOARD_ROW[(7==i ? 0 : i+1)][j], // e
                                        BOARD_ROW[(7==i ? 0 : i+1)][(0==j ? 7 : j-1)], // se
                                        BOARD_ROW[i][(0==j ? 7 : j-1)], // s
                                        BOARD_ROW[(0==i ? 7 : i-1)][(0==j ? 7 : j-1)], // sw
                                        BOARD_ROW[(0==i ? 7 : i-1)][j], // w
                                        BOARD_ROW[(0==i ? 7 : i-1)][(7==j ? 0 : j+1)] // nw
                                       );
           end

        end

// Do these, regardless whether we are in the interactive input mode
// or running the world:

      // Sum the population total from the current state.
//    if(syncdelay[time2sum_the_rows]) // Do it always.
//      begin
         for(i=0; i<8; i=i+1) rs[i] <= c8b(BOARD_ROW[i]);
//      end

      // And compute the velocities:
      if(syncdelay[time2comp_velocities])
        begin
         for(i=0; i<8; i=i+1) 
          if(note_velocity_summed) rv[i] <= (rs[i]<<4) - (|rs[i]);
          else rv[i] <= BOARD_ROW[i][6:0];
        end

      popula <= {3'b000,rs[0]} + {3'b000,rs[1]} + {3'b000,rs[2]} + {3'b000,rs[3]}
              + {3'b000,rs[4]} + {3'b000,rs[5]} + {3'b000,rs[6]} + {3'b000,rs[7]};

//  end
  end

endmodule

